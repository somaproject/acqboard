library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


library UNISIM;
use UNISIM.VComponents.all;


-- HSEL.VHD --------------------------------------------------
-- This source generates the 18-bit twos-complement fixed-point
-- filter coefficients h[n]. Keep in mind that the output will
-- always lag one tick behind CLR due to the sync. nature of the
-- counter reset and sync nature of the ram.  
entity HSEL is
    Port ( CLK2X : in std_logic;
           CLR : in std_logic;
			  RESET : in std_logic; 
           HD : out std_logic_vector(21 downto 0));
end HSEL;

architecture Behavioral of HSEL is
	signal index: std_logic_vector(7 downto 0) := "00000000"; 
	signal hdl: std_logic_vector(21 downto 0); 		  

	signal DO_Dummy: std_logic_vector(9 downto 0); 
	component RAMB4_S16
		generic (
	       INIT_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000");
	  port (DI     : in STD_LOGIC_VECTOR (15 downto 0);
	        EN     : in STD_logic;
	        WE     : in STD_logic;
	        RST    : in STD_logic;
	        CLK    : in STD_logic;
	        ADDR   : in STD_LOGIC_VECTOR (7 downto 0);
	        DO     : out STD_LOGIC_VECTOR (15 downto 0)); 
	end component;

begin
	
	-- counter vhdl
	counter: process(CLK2X) is
	begin
		if rising_edge(CLK2X) then
			if CLR = '1' then
				index <= "00000000";
				--HD <= "0000000000000000000000";
			else
				index <= index + 1;
				--HD <= hdl;
			end if;
		end if; 
	
	end process counter;  
	HD <= hdl; 
	-- RAM instantiation

	RAML: RAMB4_S16 
		generic map (
			INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
			)
		port map (
			DI =>	"0000000000000000",
			EN => '1',
			WE => '0',
			RST => CLR,
			CLK => CLK2X,
			ADDR => 	index,
			DO => hdl(15 downto 0));

	RAMH: RAMB4_S16 
		generic map (
			INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000020",
			INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
			)
		port map (
			DI =>	"0000000000000000",
			EN => '1',
			WE => '0',
			RST => CLR,
			CLK => CLK2X,
			ADDR => 	index,
			DO(5 downto 0) => hdl(21 downto 16),
			DO(15 downto 6)  => DO_dummy);


end Behavioral;
