library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


library UNISIM;
use UNISIM.VComponents.all;


-- HSEL.VHD --------------------------------------------------
-- This source generates the 18-bit twos-complement fixed-point
-- filter coefficients h[n]. Keep in mind that the output will
-- always lag one tick behind CLR due to the sync. nature of the
-- counter reset and sync nature of the ram.  
entity HSEL is
    Port ( CLK2X : in std_logic;
           CLR : in std_logic;
			  RESET : in std_logic; 
           HD : out std_logic_vector(21 downto 0));
end HSEL;

architecture Behavioral of HSEL is
	signal index: std_logic_vector(7 downto 0) := "00000000"; 
	signal hdl: std_logic_vector(21 downto 0); 		  

	signal DO_Dummy: std_logic_vector(9 downto 0); 
	component RAMB4_S16
		generic (
	       INIT_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000");
	  port (DI     : in STD_LOGIC_VECTOR (15 downto 0);
	        EN     : in STD_logic;
	        WE     : in STD_logic;
	        RST    : in STD_logic;
	        CLK    : in STD_logic;
	        ADDR   : in STD_LOGIC_VECTOR (7 downto 0);
	        DO     : out STD_LOGIC_VECTOR (15 downto 0)); 
	end component;

begin
	
	-- counter vhdl
	counter: process(CLK2X) is
	begin
		if rising_edge(CLK2X) then
			if CLR = '1' then
				index <= "00000000";
				HD <= "0000000000000000000000";
			else
				index <= index + 1;
				HD <= hdl;
			end if;
		end if; 
	
	end process counter;  
	
	-- RAM instantiation

	RAML: RAMB4_S16 
		generic map (
			--INIT_00 => X"EDA4F15AF4DDF803FAAEFCD4FE73FF96005000B300D700D100B10086005A0049",
			--INIT_01 => X"379C318328B01E1812B1075BFCD3F3AEEC50E6EFE394E223E261E400E6A7E9FA",
			--INIT_02 => X"B4E394DA81A37A757DEE8A3D9D41B4B7CE5FE821002C150925AB317538343A16",
			--INIT_03 => X"7ADAA779C32BCC8EC32BA7797ADA3F7FF84CA8A35437FECCAC065F311B15E1D8",
			--INIT_04 => X"9D418A3D7DEE7A7581A394DAB4E3E1D81B155F31AC06FECC5437A8A3F84C3F7F",
			--INIT_05 => X"FCD3075B12B11E1828B03183379C3A163834317525AB1509002CE821CE5FB4B7",
			--INIT_06 => X"FE73FCD4FAAEF803F4DDF15AEDA4E9FAE6A7E400E261E223E394E6EFEC50F3AE",
			--INIT_07 => X"00000000000000000000000000000049005A008600B100D100D700B30050FF96"
			)
		port map (
			DI =>	"0000000000000000",
			EN => '1',
			WE => '0',
			RST => CLR,
			CLK => CLK2X,
			ADDR => 	index,
			DO => hdl(15 downto 0));

	RAMH: RAMB4_S16 
		generic map (
			--INIT_00 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000",
			--INIT_01 => X"000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
			--INIT_02 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000",
			--INIT_03 => X"000200020002000200020002000200020001000100010000000000000000FFFF",
			--INIT_04 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000001000100010002",
			--INIT_05 => X"FFFF000000000000000000000000000000000000000000000000FFFFFFFFFFFF",
			--INIT_06 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
			--INIT_07 => X"000000000000000000000000000000000000000000000000000000000000FFFF"
			)
		port map (
			DI =>	"0000000000000000",
			EN => '1',
			WE => '0',
			RST => CLR,
			CLK => CLK2X,
			ADDR => 	index,
			DO(5 downto 0) => hdl(21 downto 16),
			DO(15 downto 6)  => DO_dummy);


end Behavioral;
